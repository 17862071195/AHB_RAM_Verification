`ifndef AHB_RAM_TESTS_SVH
`define AHB_RAM_TESTS_SVH

`include "ahb_ram_base_test.sv"
`include "ahb_ram_smoke_test.sv"
`include "ahb_ram_diff_hsize_test.sv"
`include "ahb_ram_diff_haddr_test.sv"
`include "ahb_ram_reset_w2r_test.sv"
`include "ahb_ram_haddr_word_unaligned_test.sv"

`endif // AHB_RAM_TESTS_SVH
