`ifndef AHB_RAM_PKG_SV
`define AHB_RAM_PKG_SV

package ahb_ram_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import lvc_ahb_pkg::*;

  `include "ahb_ram_reg.sv"
  `include "ahb_ram_reg_adapter.sv"
  `include "ahb_ram_config.sv"
  `include "ahb_ram_subscriber.sv"
  `include "ahb_ram_scoreboard.sv"
  `include "ahb_ram_cov.sv"
  `include "ahb_ram_virtual_sequencer.sv"
  `include "ahb_ram_env.sv"
  `include "ahb_ram_seq_lib.svh"
  `include "ahb_ram_tests.svh"

  
endpackage

`endif //AHB_RAM_PKG_SV
