`ifndef AHB_RAM_ELEMENT_SEQUENCES_SVH
`define AHB_RAM_ELEMENT_SEQUENCES_SVH

  `include "ahb_ram_base_element_sequence.sv"
  `include "ahb_ram_single_write_seq.sv"
  `include "ahb_ram_single_read_seq.sv"

`endif // AHB_RAM_ELEMENT_SEQUENCES_SVH
