`ifndef AHB_RAM_TESTS_SVH
`define AHB_RAM_TESTS_SVH

`include "ahb_ram_base_test.sv"
`include "ahb_ram_smoke_test.sv"

`endif // AHB_RAM_TESTS_SVH
