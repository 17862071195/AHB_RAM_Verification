`ifndef AHB_RAM_SEQ_LIB_SVH
`define AHB_RAM_SEQ_LIB_SVH

`include "ahb_ram_element_sequences.svh"
`include "ahb_ram_base_virtual_sequence.sv"
`include "ahb_ram_smoke_virt_seq.sv"
`include "ahb_ram_diff_hsize_virt_seq.sv"
`include "ahb_ram_diff_haddr_virt_seq.sv"

`endif // AHB_RAM_SEQ_LIB_SVH
