`ifndef AHB_RAM_SEQ_LIB_SVH
`define AHB_RAM_SEQ_LIB_SVH

`include "ahb_ram_base_virtual_sequence.sv"
`include "ahb_ram_smoke_virt_seq.sv"

`endif // AHB_RAM_SEQ_LIB_SVH
