`ifndef AHB_RAM_IF_SV
`define AHB_RAM_IF_SV

interface ahb_ram_if;
  logic clk;
  logic rstn;
  

endinterface

`endif //AHB_RAM_IF_SV

