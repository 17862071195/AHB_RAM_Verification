`ifndef LVC_AHB_IF_SV
`define LVC_AHB_IF_SV

interface lvc_ahb_if;

endinterface
`endif //LVC_AHB_IF_SV
