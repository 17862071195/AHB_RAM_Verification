`ifndef LVC_AHB_SEQUENCE_LIB_SVH
`define LVC_AHB_SEQUENCE_LIB_SVH

  `include "lvc_ahb_base_sequence.sv"
  `include "lvc_ahb_master_single_trnas.sv"

`endif // LVC_AHB_SEQUENCE_LIB_SVH
